class ALU_item;

    rand bit [3:0]  A,B;
    rand bit [1:0]  ALU_FUN;
         bit        CLK;
         bit [7:0] ALU_OUT;
endclass