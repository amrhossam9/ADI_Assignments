interface ALU_if(input bit CLK);
   logic [3:0]  A, B;
   logic [1:0]  ALU_FUN;
   logic [7:0]  ALU_OUT;
endinterface
